/////////////////////////////////////////////////////////////////////
// ---------------------- IVCAD 2018 Spring ---------------------- //
// ---------------------- Editor : JohnChang ----------------------//
// ---------------------- Date : 2018.03    ---------------------- //
// ----------------------      test1        ---------------------- // 
/////////////////////////////////////////////////////////////////////
module test1(out1, 
             out2,
             in1, 
             in2);
             
input   in1 , in2;
output  out1 , out2;
	
assign out1 = in1 & in2;	//and
assign out2 = in1 | in2;	//or
	
endmodule