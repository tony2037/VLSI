/////////////////////////////////////////////////////////////////////
// ---------------------- IVCAD 2018 Spring ---------------------- //
// ---------------------- Editor : JohnChang ----------------------//
// ---------------------- Date : 2018.03    ---------------------- //
// ----------------------      test2        ---------------------- // 
/////////////////////////////////////////////////////////////////////
module test2(out1, 
             out2,
             out3, 
             in1, 
             in2);
            
input  in1, in2;
output out1 ,out2, out3;

assign out1 = ~in2;         //not
assign out2 = in1 | in2;   //or
assign out3 = in1 ^ in2;   //xor

endmodule
